library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Priorità: Preset -> Clear -> Clock -> Data

entity LatchPCP is
    Port ( D, clk, clr, pre : in  STD_LOGIC;
           Q : out  STD_LOGIC);
end LatchPCP;

architecture Behavioral of LatchPCP is
    begin
        process(clk, D, clr, pre)
            begin
                if(pre = '1') then -- Se il Preset è attivo (1 Poichè Latch Positivo, 0 Se Negativo)
                    Q <= '1'; -- Allora assegno 1 all'uscita Q
                else if(clr = '1') then -- Se il Reset è attivo (1 Poichè Latch Positivo, 0 Se Negativo)
                    Q <= '0'; -- Allora assegno 0 all'uscita Q
                else if(clk = '1') then -- Se il Clock è attivo (1 Poichè Latch Positivo, 0 Se Negativo)
                    Q <= D; -- Allora assegno il valore d'ingresso D all'uscita Q
                end if;
        end process;
end Behavioral;